** sch_path: /home/shr25031/ihp-mpw-be/ihp-mpw-be/TO_Apr2025/Mixer5GHz/xschem/Mixer5GHz.sch
.subckt Mixer5GHz RFN RFP VDC IFP IFN IDC OSCN OSCP VCC ICC GND
*.PININFO RFN:B RFP:B VDC:B IFP:B IFN:B IDC:B OSCN:B OSCP:B VCC:B ICC:B GND:B
M6 RFN LON net2 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XRL2 RFN VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XRL1 RFP VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
M8 RFN LOP net3 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
M7 RFP LON net3 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
M5 RFP LOP net2 GND sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
M4 net3 IFN net1 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
M3 net2 IFP net1 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
M2 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
M1 net1 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
M11 LOP LON net4 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
M12 LON LOP net4 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
M9 IDC IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
M10 net4 IDC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XC1 VDC LOP cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR1 LOP VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XC2 VDC LON cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR2 LON VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
M13 OSCP OSCN net5 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
M14 OSCN OSCP net5 GND sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
M15 ICC ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
M16 net5 ICC GND GND sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XC3 VCC OSCP cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR3 OSCP VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XC4 VCC OSCN cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR4 OSCN VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XL1 VDC LOP GND inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
XL2 VDC LON GND inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
XL3 VCC OSCP GND inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
XL4 VCC OSCN GND inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
.ends
