** sch_path: /home/shr25031/ihp-mpw-be/ihp-mpw-be/TO_Apr2025/Mixer5GHz/xschem/Mixer5GHz.sch
.subckt Mixer5GHz RFN RFP VDC IFP IFN IDC OSCN OSCP VCC ICC GNDC GNDD
*.PININFO RFN:B RFP:B VDC:B IFP:B IFN:B IDC:B OSCN:B OSCP:B VCC:B ICC:B GNDC:B GNDD:B
XM6 RFN LON net2 GNDD sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XRL2 RFN VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XRL1 RFP VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XM8 RFN LOP net3 GNDD sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XM7 RFP LON net3 GNDD sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XM5 RFP LOP net2 GNDD sg13_lv_nmos w=60.0u l=0.13u ng=10 m=1
XM4 net3 IFN net1 GNDD sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM3 net2 IFP net1 GNDD sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM2 IDC IDC GNDD GNDD sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM1 net1 IDC GNDD GNDD sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM11 LOP LON net4 GNDD sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM12 LON LOP net4 GNDD sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM9 IDC IDC GNDD GNDD sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM10 net4 IDC GNDD GNDD sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XC1 VDC LOP cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR1 LOP VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XC2 VDC LON cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR2 LON VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XM13 OSCP OSCN net5 GNDC sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM14 OSCN OSCP net5 GNDC sg13_lv_nmos w=90.0u l=0.13u ng=15 m=1
XM15 ICC ICC GNDC GNDC sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XM16 net5 ICC GNDC GNDC sg13_lv_nmos w=120.0u l=0.13u ng=20 m=1
XC3 VCC OSCP cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR3 OSCP VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XC4 VCC OSCN cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR4 OSCN VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XL1 VDC LOP GNDD inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
XL2 VDC LON GNDD inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
XL3 VCC OSCP GNDC inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
XL4 VCC OSCN GNDC inductor2 w=10e-6 s=10e-6 d=222e-6 nr_r=2 m=1
.ends
