** sch_path: /home/shr25031/ihp-mpw-be/ihp-mpw-be/TO_Apr2025/160GHz_LNA/xschem/160GHz_LNA.sch
.subckt 160GHz_LNA RF_INPUT GND VCC VBB1 RF_OUTPUT VBB2
*.PININFO RF_INPUT:I GND:B VCC:B VBB1:B RF_OUTPUT:O VBB2:B
XC1 RF_INPUT net1 GND rfcmim w=10.0e-6 l=15.0e-6 wfeed=6.0e-6
XQ1 net2 net1 GND GND npn13G2 le=900e-9 we=70.0n m=4
XRc1 net2 VCC rsil w=7.5e-6 l=5.0e-6 m=1 b=0
XRb1 net1 VBB1 rhigh w=1.9e-6 l=6.0e-6 m=1 b=0
XCDecap1 VBB1 GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XCDecap2 VCC GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XC2 net2 GND GND rfcmim w=32.0e-6 l=3.72e-6 wfeed=3.0e-6
XC3 GND net3 GND rfcmim w=5.2e-6 l=2.4e-6 wfeed=3.0e-6
XRb2 net3 VBB1 rhigh w=1.9e-6 l=5.0e-6 m=1 b=0
XCDecap3 VBB1 GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XQ2 net4 net3 GND GND npn13G2 le=900e-9 we=70.0n m=4
XRc2 net4 VCC rsil w=7.5e-6 l=5.0e-6 m=1 b=0
XCDecap4 VCC GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XC4 net4 GND GND rfcmim w=32.0e-6 l=3.72e-6 wfeed=3.0e-6
XC5 GND net5 GND rfcmim w=7.6e-6 l=2.5e-6 wfeed=3.0e-6
XRb3 net5 VBB1 rhigh w=1.9e-6 l=6.0e-6 m=1 b=0
XCDecap5 VBB1 GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XRc3 net6 VCC rsil w=7.5e-6 l=5.0e-6 m=1 b=0
XCDecap6 VCC GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XQ3 net6 net5 GND GND npn13G2 le=900e-9 we=70.0n m=2
XRb4 net7 VBB2 rhigh w=2.0e-6 l=6.0e-6 m=1 b=0
XCDecap7 VBB2 GND cap_cmim w=20.0e-6 l=25.0e-6 m=4
XRc4 net8 VCC rsil w=7.5e-6 l=5.5e-6 m=1 b=0
XCDecap8 VCC GND cap_cmim w=20.0e-6 l=25.0e-6 m=2
XQ4 net8 net7 GND GND npn13G2 le=900e-9 we=70.0n m=2
XC6 net6 GND GND rfcmim w=32.0e-6 l=12.5e-6 wfeed=3.0e-6
XC7 GND net7 GND rfcmim w=5.1e-6 l=2.4e-6 wfeed=3.0e-6
XC8 net8 GND GND rfcmim w=32.0e-6 l=6.2e-6 wfeed=3.0e-6
XC9 GND RF_OUTPUT GND rfcmim w=3.2e-6 l=2.4e-6 wfeed=3.0e-6
.ends
