** sch_path: /home/shr25031/ihp-mpw-be/ihp-mpw-be/TO_Apr2025/Mixer5GHz/xschem/Mixer5GHz.sch
.subckt Mixer5GHz RFN RFP VDC IFP IFN GND IDC OSCN OSCP VCC ICC GND
*.PININFO RFN:B RFP:B VDC:B IFP:B IFN:B GND:B IDC:B OSCN:B OSCP:B VCC:B ICC:B GND:B
XM6 net2 LON RFN GND sg13_lv_nmos l=0.13u w=60.0u ng=10 m=1
XRL2 RFN VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XRL1 RFP VDC rppd w=4.50e-6 l=3.20e-6 m=1 b=0
XM8 net3 LOP RFN GND sg13_lv_nmos l=0.13u w=60.0u ng=10 m=1
XM7 net3 LON RFP GND sg13_lv_nmos l=0.13u w=60.0u ng=10 m=1
XM5 net2 LOP RFP GND sg13_lv_nmos l=0.13u w=60.0u ng=10 m=1
XM4 net1 IFN net3 GND sg13_lv_nmos l=0.13u w=90.0u ng=15 m=1
XM3 net1 IFP net2 GND sg13_lv_nmos l=0.13u w=90.0u ng=15 m=1
XM2 GND IDC IDC GND sg13_lv_nmos l=0.13u w=120.0u ng=20 m=1
XM1 GND IDC net1 GND sg13_lv_nmos l=0.13u w=120.0u ng=20 m=1
XM11 net4 LON LOP GND sg13_lv_nmos l=0.13u w=90.0u ng=15 m=1
XM12 net4 LOP LON GND sg13_lv_nmos l=0.13u w=90.0u ng=15 m=1
XM9 GND IDC IDC GND sg13_lv_nmos l=0.13u w=120.0u ng=20 m=1
XM10 GND IDC net4 GND sg13_lv_nmos l=0.13u w=120.0u ng=20 m=1
XC1 VDC LOP cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR1 LOP VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XC2 VDC LON cap_cmim w=11.745e-6 l=9.445e-6 m=1
XR2 LON VDC rppd w=4.4e-6 l=1.5e-6 m=1 b=0
XM13 net5 OSCN OSCP GND sg13_lv_nmos l=0.13u w=90.0u ng=15 m=1
XM14 net5 OSCP OSCN GND sg13_lv_nmos l=0.13u w=90.0u ng=15 m=1
XM15 GND ICC ICC GND sg13_lv_nmos l=0.13u w=120.0u ng=20 m=1
XM16 GND ICC net5 GND sg13_lv_nmos l=0.13u w=120.0u ng=20 m=1
XC3 VCC OSCP cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR3 OSCP VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
XC4 VCC OSCN cap_cmim w=19.1e-6 l=10.7e-6 m=1
XR4 OSCN VCC rppd w=4.35e-6 l=1.5e-6 m=1 b=0
L3 VCC OSCP 2.006n m=1
L1 VDC LOP 2.006n m=1
L2 VDC LON 2.006n m=1
L4 VCC OSCN 2.006n m=1
.ends
